VERSION 5.7 ;
BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.17 ;
END li1

LAYER mcon
  TYPE CUT ;
END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.34 ;
  WIDTH 0.14 ;
END met1

LAYER via
  TYPE CUT ;
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.46 ;
  WIDTH 0.14 ;
END met2

LAYER via2
  TYPE CUT ;
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.68 ;
  WIDTH 0.3 ;
END met3

LAYER via3
  TYPE CUT ;
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.92 ;
  WIDTH 0.3 ;
END met4

LAYER via4
  TYPE CUT ;
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3.4 ;
  WIDTH 1.6 ;
END met5

LAYER nwell
  TYPE MASTERSLICE ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
END pwell

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA L1M1_PR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C
  LAYER li1 ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER mcon ;
    RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
    RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_Enc

VIA M1M2_PR_R
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_R_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_R_Enc

VIA M1M2_PR_M
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_M_Enc
  LAYER met1 ;
    RECT -0.16 -0.13 0.16 0.13 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_M_Enc

VIA M1M2_PR_MR
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_MR_Enc
  LAYER met1 ;
    RECT -0.13 -0.16 0.13 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_MR_Enc

VIA M1M2_PR_C
  LAYER met1 ;
    RECT -0.16 -0.16 0.16 0.16 ;
  LAYER via ;
    RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met2 ;
    RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M
  LAYER met2 ;
    RECT -0.14 -0.185 0.14 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR
  LAYER met2 ;
    RECT -0.185 -0.14 0.185 0.14 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C
  LAYER met2 ;
    RECT -0.185 -0.185 0.185 0.185 ;
  LAYER via2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M
  LAYER met3 ;
    RECT -0.19 -0.16 0.19 0.16 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR
  LAYER met3 ;
    RECT -0.16 -0.19 0.16 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C
  LAYER met3 ;
    RECT -0.19 -0.19 0.19 0.19 ;
  LAYER via3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met4 ;
    RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C
  LAYER met4 ;
    RECT -0.59 -0.59 0.59 0.59 ;
  LAYER via4 ;
    RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met5 ;
    RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

SITE unit
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.46 BY 2.72 ;
END unit

SITE unithddbl
  CLASS CORE ;
  SIZE 0.46 BY 5.44 ;
END unithddbl

MACRO sb_1__0_
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 139.84 BY 103.36 ;
  SYMMETRY X Y ;
  PIN pReset[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.96 102 60.1 103.36 ;
    END
  END pReset[0]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.62 102 69.76 103.36 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.04 102 36.18 103.36 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.23 102 93.53 103.36 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.76 102 73.9 103.36 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.8 102 84.94 103.36 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.22 102 97.36 103.36 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.16 102 92.3 103.36 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.95 102 62.25 103.36 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.39 102 45.69 103.36 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.88 102 61.02 103.36 ;
    END
  END chany_top_in[9]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.83 102 75.13 103.36 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.3 102 73.44 103.36 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.06 102 53.2 103.36 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.19 102 59.49 103.36 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.96 102 106.1 103.36 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.84 102 95.98 103.36 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.6 102 98.74 103.36 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.4 102 89.54 103.36 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.27 102 81.57 103.36 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.66 102 34.8 103.36 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.04 102 59.18 103.36 ;
    END
  END chany_top_in[20]
  PIN chany_top_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.94 102 43.08 103.36 ;
    END
  END chany_top_in[21]
  PIN chany_top_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.42 102 83.56 103.36 ;
    END
  END chany_top_in[22]
  PIN chany_top_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.03 102 84.33 103.36 ;
    END
  END chany_top_in[23]
  PIN chany_top_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 98.75 102 99.05 103.36 ;
    END
  END chany_top_in[24]
  PIN chany_top_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.99 102 96.29 103.36 ;
    END
  END chany_top_in[25]
  PIN chany_top_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.84 102 72.98 103.36 ;
    END
  END chany_top_in[26]
  PIN chany_top_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.18 102 86.32 103.36 ;
    END
  END chany_top_in[27]
  PIN chany_top_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.98 102 100.12 103.36 ;
    END
  END chany_top_in[28]
  PIN chany_top_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.56 102 87.7 103.36 ;
    END
  END chany_top_in[29]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 31.28 96.07 32.66 96.37 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_[0]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.32 85.68 21.46 87.04 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_[0]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.96 85.68 14.1 87.04 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_[0]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.1 85.68 18.24 87.04 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_[0]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 31.28 96.32 31.875 96.46 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_[0]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.18 85.68 17.32 87.04 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_[0]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 31.28 97 31.875 97.14 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_[0]
  PIN top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.26 85.68 16.4 87.04 ;
    END
  END top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_[0]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 25.94 139.84 26.08 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 64.79 139.84 65.09 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 50.51 139.84 50.81 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 58.67 139.84 58.97 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 9.03 139.84 9.33 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 38.27 139.84 38.57 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 15.15 139.84 15.45 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 46.43 139.84 46.73 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 44.39 139.84 44.69 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 6.9 139.84 7.04 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 27.39 139.84 27.69 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 4.18 139.84 4.32 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 17.19 139.84 17.49 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 12.34 139.84 12.48 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 58.24 139.84 58.38 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 6.99 139.84 7.29 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 19.23 139.84 19.53 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 42.35 139.84 42.65 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 20.5 139.84 20.64 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 34.1 139.84 34.24 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 23.22 139.84 23.36 ;
    END
  END chanx_right_in[20]
  PIN chanx_right_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 33.51 139.84 33.81 ;
    END
  END chanx_right_in[21]
  PIN chanx_right_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 77.03 139.84 77.33 ;
    END
  END chanx_right_in[22]
  PIN chanx_right_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 72.95 139.84 73.25 ;
    END
  END chanx_right_in[23]
  PIN chanx_right_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 15.06 139.84 15.2 ;
    END
  END chanx_right_in[24]
  PIN chanx_right_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 56.63 139.84 56.93 ;
    END
  END chanx_right_in[25]
  PIN chanx_right_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 55.86 139.84 56 ;
    END
  END chanx_right_in[26]
  PIN chanx_right_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 74.99 139.84 75.29 ;
    END
  END chanx_right_in[27]
  PIN chanx_right_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 17.44 139.84 17.58 ;
    END
  END chanx_right_in[28]
  PIN chanx_right_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 80 139.84 80.14 ;
    END
  END chanx_right_in[29]
  PIN right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 14.38 139.84 14.52 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 33.42 139.84 33.56 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 4.95 139.84 5.25 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 80.68 139.84 80.82 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 3.59 139.84 3.89 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 1.8 139.84 1.94 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 77.96 139.84 78.1 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 36.23 139.84 36.53 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_[0]
  PIN right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 75.24 139.84 75.38 ;
    END
  END right_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_[0]
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 6.9 0.595 7.04 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 69.55 1.38 69.85 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 20.5 0.595 20.64 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 69.12 0.595 69.26 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 82.47 1.38 82.77 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 25.35 1.38 25.65 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 9.62 0.595 9.76 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 38.27 1.38 38.57 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 19.23 1.38 19.53 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 23.31 1.38 23.61 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 33.51 1.38 33.81 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 13.11 1.38 13.41 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 31.47 1.38 31.77 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 60.96 0.595 61.1 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 66.4 0.595 66.54 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 55.86 0.595 56 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 62.75 1.38 63.05 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 80.43 1.38 80.73 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 15.06 0.595 15.2 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 71.84 0.595 71.98 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 15.15 1.38 15.45 ;
    END
  END chanx_left_in[20]
  PIN chanx_left_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 75.67 1.38 75.97 ;
    END
  END chanx_left_in[21]
  PIN chanx_left_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 63.68 0.595 63.82 ;
    END
  END chanx_left_in[22]
  PIN chanx_left_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 73.63 1.38 73.93 ;
    END
  END chanx_left_in[23]
  PIN chanx_left_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 44.39 1.38 44.69 ;
    END
  END chanx_left_in[24]
  PIN chanx_left_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 77.28 0.595 77.42 ;
    END
  END chanx_left_in[25]
  PIN chanx_left_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 71.59 1.38 71.89 ;
    END
  END chanx_left_in[26]
  PIN chanx_left_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 46.43 1.38 46.73 ;
    END
  END chanx_left_in[27]
  PIN chanx_left_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 60.71 1.38 61.01 ;
    END
  END chanx_left_in[28]
  PIN chanx_left_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 21.27 1.38 21.57 ;
    END
  END chanx_left_in[29]
  PIN left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 17.44 0.595 17.58 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 4.27 1.38 4.57 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 9.71 1.38 10.01 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 77.71 1.38 78.01 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 8.35 1.38 8.65 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 1.8 0.595 1.94 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 6.99 1.38 7.29 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 55.18 0.595 55.32 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_[0]
  PIN left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.14 0.595 36.28 ;
    END
  END left_bottom_grid_top_width_0_height_0_subtile_8__pin_inpad_0_[0]
  PIN ccff_head[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 36.14 139.84 36.28 ;
    END
  END ccff_head[0]
  PIN chany_top_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.14 102 75.28 103.36 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.94 102 66.08 103.36 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.32 102 67.46 103.36 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.32 102 44.46 103.36 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.56 102 64.7 103.36 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.06 102 76.2 103.36 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.46 102 94.6 103.36 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.51 102 78.81 103.36 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.04 102 82.18 103.36 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.82 102 78.96 103.36 ;
    END
  END chany_top_out[9]
  PIN chany_top_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.8 102 38.94 103.36 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.28 102 56.42 103.36 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.68 102 74.82 103.36 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.54 102 70.68 103.36 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.38 102 49.52 103.36 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.78 102 90.92 103.36 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.26 102 62.4 103.36 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.22 102 74.36 103.36 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.44 102 77.58 103.36 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.15 102 48.45 103.36 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.11 102 37.41 103.36 ;
    END
  END chany_top_out[20]
  PIN chany_top_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.58 102 104.72 103.36 ;
    END
  END chany_top_out[21]
  PIN chany_top_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.44 102 54.58 103.36 ;
    END
  END chany_top_out[22]
  PIN chany_top_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.08 102 47.22 103.36 ;
    END
  END chany_top_out[23]
  PIN chany_top_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.47 102 90.77 103.36 ;
    END
  END chany_top_out[24]
  PIN chany_top_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.7 102 68.84 103.36 ;
    END
  END chany_top_out[25]
  PIN chany_top_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.42 102 37.56 103.36 ;
    END
  END chany_top_out[26]
  PIN chany_top_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.08 102 70.22 103.36 ;
    END
  END chany_top_out[27]
  PIN chany_top_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.76 102 50.9 103.36 ;
    END
  END chany_top_out[28]
  PIN chany_top_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.66 102 80.8 103.36 ;
    END
  END chany_top_out[29]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 74.56 139.84 74.7 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 80.43 139.84 80.73 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 40.31 139.84 40.61 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 77.28 139.84 77.42 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 31.04 139.84 31.18 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 9.62 139.84 9.76 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 39.2 139.84 39.34 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 71.84 139.84 71.98 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 69.12 139.84 69.26 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 50.42 139.84 50.56 ;
    END
  END chanx_right_out[9]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 41.92 139.84 42.06 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 82.72 139.84 82.86 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 36.82 139.84 36.96 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 13.11 139.84 13.41 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 82.47 139.84 82.77 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 64.02 139.84 64.16 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 52.55 139.84 52.85 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 47.7 139.84 47.84 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 44.64 139.84 44.78 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 68.87 139.84 69.17 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 53.14 139.84 53.28 ;
    END
  END chanx_right_out[20]
  PIN chanx_right_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 66.4 139.84 66.54 ;
    END
  END chanx_right_out[21]
  PIN chanx_right_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 31.47 139.84 31.77 ;
    END
  END chanx_right_out[22]
  PIN chanx_right_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 70.91 139.84 71.21 ;
    END
  END chanx_right_out[23]
  PIN chanx_right_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 29.43 139.84 29.73 ;
    END
  END chanx_right_out[24]
  PIN chanx_right_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 61.39 139.84 61.69 ;
    END
  END chanx_right_out[25]
  PIN chanx_right_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 60.96 139.84 61.1 ;
    END
  END chanx_right_out[26]
  PIN chanx_right_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 48.47 139.84 48.77 ;
    END
  END chanx_right_out[27]
  PIN chanx_right_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 28.66 139.84 28.8 ;
    END
  END chanx_right_out[28]
  PIN chanx_right_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 66.83 139.84 67.13 ;
    END
  END chanx_right_out[29]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 40.31 1.38 40.61 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 52.8 0.595 52.94 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 29.43 1.38 29.73 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 12.34 0.595 12.48 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 42.35 1.38 42.65 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 17.19 1.38 17.49 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 31.38 0.595 31.52 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 50.42 0.595 50.56 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 4.18 0.595 4.32 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 47.7 0.595 47.84 ;
    END
  END chanx_left_out[9]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 41.92 0.595 42.06 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 80 0.595 80.14 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 25.94 0.595 26.08 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 74.56 0.595 74.7 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 27.39 1.38 27.69 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 58.24 0.595 58.38 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 39.2 0.595 39.34 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 50.51 1.38 50.81 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 23.22 0.595 23.36 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 82.72 0.595 82.86 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 48.47 1.38 48.77 ;
    END
  END chanx_left_out[20]
  PIN chanx_left_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 58.67 1.38 58.97 ;
    END
  END chanx_left_out[21]
  PIN chanx_left_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 36.82 0.595 36.96 ;
    END
  END chanx_left_out[22]
  PIN chanx_left_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 67.51 1.38 67.81 ;
    END
  END chanx_left_out[23]
  PIN chanx_left_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 28.66 0.595 28.8 ;
    END
  END chanx_left_out[24]
  PIN chanx_left_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 56.63 1.38 56.93 ;
    END
  END chanx_left_out[25]
  PIN chanx_left_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 44.64 0.595 44.78 ;
    END
  END chanx_left_out[26]
  PIN chanx_left_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 52.55 1.38 52.85 ;
    END
  END chanx_left_out[27]
  PIN chanx_left_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 34.1 0.595 34.24 ;
    END
  END chanx_left_out[28]
  PIN chanx_left_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 64.79 1.38 65.09 ;
    END
  END chanx_left_out[29]
  PIN ccff_tail[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 5.63 1.38 5.93 ;
    END
  END ccff_tail[0]
  PIN pReset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.8 0 61.94 1.36 ;
    END
  END pReset_S_in
  PIN pReset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.66 102 57.8 103.36 ;
    END
  END pReset_N_out
  PIN pReset_W_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0 36.23 1.38 36.53 ;
    END
  END pReset_W_out
  PIN pReset_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 139.245 85.1 139.84 85.24 ;
    END
  END pReset_E_out
  PIN Test_en_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.4 0 66.54 1.36 ;
    END
  END Test_en_S_in
  PIN Test_en_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.7 102 45.84 103.36 ;
    END
  END Test_en_N_out
  PIN reset_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.72 0 62.86 1.36 ;
    END
  END reset_S_in
  PIN reset_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.36 102 101.5 103.36 ;
    END
  END reset_N_out
  PIN sc_head_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0 18.12 0.595 18.26 ;
    END
  END sc_head_W_in
  PIN sc_head_E_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.46 21.27 139.84 21.57 ;
    END
  END sc_head_E_out
  PIN prog_clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met2 ;
        RECT 63.64 102 63.78 103.36 ;
    END
  END prog_clk
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER met4 ;
        RECT 51.83 102 52.13 103.36 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_1_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.75 0 76.05 1.36 ;
    END
  END prog_clk_1_S_in
  PIN prog_clk_1_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 65.63 102 65.93 103.36 ;
    END
  END prog_clk_1_N_out
  PIN clk_2_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.31 0 69.61 0.8 ;
    END
  END clk_2_S_in
  PIN clk_2_N_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.31 102.56 69.61 103.36 ;
    END
  END clk_2_N_out
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 0 10.52 4.8 15.32 ;
        RECT 135.04 10.52 139.84 15.32 ;
        RECT 0 54.52 4.8 59.32 ;
        RECT 135.04 54.52 139.84 59.32 ;
      LAYER met4 ;
        RECT 19.33 0 20.83 1.5 ;
        RECT 39.73 0 41.23 1.5 ;
        RECT 70.97 0 72.47 1.5 ;
        RECT 102.21 0 103.71 1.5 ;
        RECT 126.21 0 127.71 1.5 ;
        RECT 19.33 85.54 20.83 87.04 ;
        RECT 126.21 85.54 127.71 87.04 ;
        RECT 39.73 101.86 41.23 103.36 ;
        RECT 70.97 101.86 72.47 103.36 ;
        RECT 102.21 101.86 103.71 103.36 ;
      LAYER met1 ;
        RECT 0 -0.24 0.48 0.24 ;
        RECT 139.36 -0.24 139.84 0.24 ;
        RECT 0 5.2 0.48 5.68 ;
        RECT 139.36 5.2 139.84 5.68 ;
        RECT 0 10.64 0.48 11.12 ;
        RECT 139.36 10.64 139.84 11.12 ;
        RECT 0 16.08 0.48 16.56 ;
        RECT 139.36 16.08 139.84 16.56 ;
        RECT 0 21.52 0.48 22 ;
        RECT 139.36 21.52 139.84 22 ;
        RECT 0 26.96 0.48 27.44 ;
        RECT 139.36 26.96 139.84 27.44 ;
        RECT 0 32.4 0.48 32.88 ;
        RECT 139.36 32.4 139.84 32.88 ;
        RECT 0 37.84 0.48 38.32 ;
        RECT 139.36 37.84 139.84 38.32 ;
        RECT 0 43.28 0.48 43.76 ;
        RECT 139.36 43.28 139.84 43.76 ;
        RECT 0 48.72 0.48 49.2 ;
        RECT 139.36 48.72 139.84 49.2 ;
        RECT 0 54.16 0.48 54.64 ;
        RECT 139.36 54.16 139.84 54.64 ;
        RECT 0 59.6 0.48 60.08 ;
        RECT 139.36 59.6 139.84 60.08 ;
        RECT 0 65.04 0.48 65.52 ;
        RECT 139.36 65.04 139.84 65.52 ;
        RECT 0 70.48 0.48 70.96 ;
        RECT 139.36 70.48 139.84 70.96 ;
        RECT 0 75.92 0.48 76.4 ;
        RECT 139.36 75.92 139.84 76.4 ;
        RECT 0 81.36 0.48 81.84 ;
        RECT 139.36 81.36 139.84 81.84 ;
        RECT 0 86.8 0.48 87.28 ;
        RECT 139.36 86.8 139.84 87.28 ;
        RECT 31.28 92.24 31.76 92.72 ;
        RECT 108.08 92.24 108.56 92.72 ;
        RECT 31.28 97.68 31.76 98.16 ;
        RECT 108.08 97.68 108.56 98.16 ;
        RECT 31.28 103.12 31.76 103.6 ;
        RECT 108.08 103.12 108.56 103.6 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0 32.52 4.8 37.32 ;
        RECT 135.04 32.52 139.84 37.32 ;
        RECT 0 76.52 4.8 81.32 ;
        RECT 135.04 76.52 139.84 81.32 ;
      LAYER met4 ;
        RECT 3.71 0 5.21 1.5 ;
        RECT 55.35 0 56.85 1.5 ;
        RECT 86.59 0 88.09 1.5 ;
        RECT 3.71 85.54 5.21 87.04 ;
        RECT 55.35 101.86 56.85 103.36 ;
        RECT 86.59 101.86 88.09 103.36 ;
      LAYER met1 ;
        RECT 0 2.48 0.48 2.96 ;
        RECT 139.36 2.48 139.84 2.96 ;
        RECT 0 7.92 0.48 8.4 ;
        RECT 139.36 7.92 139.84 8.4 ;
        RECT 0 13.36 0.48 13.84 ;
        RECT 139.36 13.36 139.84 13.84 ;
        RECT 0 18.8 0.48 19.28 ;
        RECT 139.36 18.8 139.84 19.28 ;
        RECT 0 24.24 0.48 24.72 ;
        RECT 139.36 24.24 139.84 24.72 ;
        RECT 0 29.68 0.48 30.16 ;
        RECT 139.36 29.68 139.84 30.16 ;
        RECT 0 35.12 0.48 35.6 ;
        RECT 139.36 35.12 139.84 35.6 ;
        RECT 0 40.56 0.48 41.04 ;
        RECT 139.36 40.56 139.84 41.04 ;
        RECT 0 46 0.48 46.48 ;
        RECT 139.36 46 139.84 46.48 ;
        RECT 0 51.44 0.48 51.92 ;
        RECT 139.36 51.44 139.84 51.92 ;
        RECT 0 56.88 0.48 57.36 ;
        RECT 139.36 56.88 139.84 57.36 ;
        RECT 0 62.32 0.48 62.8 ;
        RECT 139.36 62.32 139.84 62.8 ;
        RECT 0 67.76 0.48 68.24 ;
        RECT 139.36 67.76 139.84 68.24 ;
        RECT 0 73.2 0.48 73.68 ;
        RECT 139.36 73.2 139.84 73.68 ;
        RECT 0 78.64 0.48 79.12 ;
        RECT 139.36 78.64 139.84 79.12 ;
        RECT 0 84.08 0.48 84.56 ;
        RECT 139.36 84.08 139.84 84.56 ;
        RECT 31.28 89.52 31.76 90 ;
        RECT 108.08 89.52 108.56 90 ;
        RECT 31.28 94.96 31.76 95.44 ;
        RECT 108.08 94.96 108.56 95.44 ;
        RECT 31.28 100.4 31.76 100.88 ;
        RECT 108.08 100.4 108.56 100.88 ;
    END
  END vssd1
  OBS
    LAYER met2 ;
      POLYGON 103.5 103.425 103.5 103.4 103.57 103.4 103.57 103.08 103.5 103.08 103.5 103.055 102.42 103.055 102.42 103.08 102.35 103.08 102.35 103.4 102.42 103.4 102.42 103.425 ;
      POLYGON 72.26 103.425 72.26 103.4 72.33 103.4 72.33 103.08 72.26 103.08 72.26 103.055 71.18 103.055 71.18 103.08 71.11 103.08 71.11 103.4 71.18 103.4 71.18 103.425 ;
      POLYGON 41.02 103.425 41.02 103.4 41.09 103.4 41.09 103.08 41.02 103.08 41.02 103.055 39.94 103.055 39.94 103.08 39.87 103.08 39.87 103.4 39.94 103.4 39.94 103.425 ;
      POLYGON 77.28 102.68 77.28 98.38 77.14 98.38 77.14 102.54 76.68 102.54 76.68 102.68 ;
      RECT 72.48 101.43 72.74 101.75 ;
      POLYGON 127.5 87.105 127.5 87.08 127.57 87.08 127.57 86.76 127.5 86.76 127.5 86.735 126.42 86.735 126.42 86.76 126.35 86.76 126.35 87.08 126.42 87.08 126.42 87.105 ;
      POLYGON 20.62 87.105 20.62 87.08 20.69 87.08 20.69 86.76 20.62 86.76 20.62 86.735 19.54 86.735 19.54 86.76 19.47 86.76 19.47 87.08 19.54 87.08 19.54 87.105 ;
      RECT 139.46 78.695 139.74 79.065 ;
      RECT 0.1 78.695 0.38 79.065 ;
      RECT 139.46 54.395 139.74 54.765 ;
      RECT 0.1 54.395 0.38 54.765 ;
      RECT 139.46 35.175 139.74 35.545 ;
      RECT 0.1 35.175 0.38 35.545 ;
      RECT 139.46 10.695 139.74 11.065 ;
      RECT 0.1 10.695 0.38 11.065 ;
      POLYGON 127.5 0.305 127.5 0.28 127.57 0.28 127.57 -0.04 127.5 -0.04 127.5 -0.065 126.42 -0.065 126.42 -0.04 126.35 -0.04 126.35 0.28 126.42 0.28 126.42 0.305 ;
      POLYGON 103.5 0.305 103.5 0.28 103.57 0.28 103.57 -0.04 103.5 -0.04 103.5 -0.065 102.42 -0.065 102.42 -0.04 102.35 -0.04 102.35 0.28 102.42 0.28 102.42 0.305 ;
      POLYGON 72.26 0.305 72.26 0.28 72.33 0.28 72.33 -0.04 72.26 -0.04 72.26 -0.065 71.18 -0.065 71.18 -0.04 71.11 -0.04 71.11 0.28 71.18 0.28 71.18 0.305 ;
      POLYGON 41.02 0.305 41.02 0.28 41.09 0.28 41.09 -0.04 41.02 -0.04 41.02 -0.065 39.94 -0.065 39.94 -0.04 39.87 -0.04 39.87 0.28 39.94 0.28 39.94 0.305 ;
      POLYGON 20.62 0.305 20.62 0.28 20.69 0.28 20.69 -0.04 20.62 -0.04 20.62 -0.065 19.54 -0.065 19.54 -0.04 19.47 -0.04 19.47 0.28 19.54 0.28 19.54 0.305 ;
      POLYGON 108.28 103.08 108.28 86.76 139.56 86.76 139.56 0.28 66.82 0.28 66.82 1.64 66.12 1.64 66.12 0.28 63.14 0.28 63.14 1.64 62.44 1.64 62.44 0.28 62.22 0.28 62.22 1.64 61.52 1.64 61.52 0.28 0.28 0.28 0.28 86.76 13.68 86.76 13.68 85.4 14.38 85.4 14.38 86.76 15.98 86.76 15.98 85.4 16.68 85.4 16.68 86.76 16.9 86.76 16.9 85.4 17.6 85.4 17.6 86.76 17.82 86.76 17.82 85.4 18.52 85.4 18.52 86.76 21.04 86.76 21.04 85.4 21.74 85.4 21.74 86.76 31.56 86.76 31.56 103.08 34.38 103.08 34.38 101.72 35.08 101.72 35.08 103.08 35.76 103.08 35.76 101.72 36.46 101.72 36.46 103.08 37.14 103.08 37.14 101.72 37.84 101.72 37.84 103.08 38.52 103.08 38.52 101.72 39.22 101.72 39.22 103.08 42.66 103.08 42.66 101.72 43.36 101.72 43.36 103.08 44.04 103.08 44.04 101.72 44.74 101.72 44.74 103.08 45.42 103.08 45.42 101.72 46.12 101.72 46.12 103.08 46.8 103.08 46.8 101.72 47.5 101.72 47.5 103.08 49.1 103.08 49.1 101.72 49.8 101.72 49.8 103.08 50.48 103.08 50.48 101.72 51.18 101.72 51.18 103.08 52.78 103.08 52.78 101.72 53.48 101.72 53.48 103.08 54.16 103.08 54.16 101.72 54.86 101.72 54.86 103.08 56 103.08 56 101.72 56.7 101.72 56.7 103.08 57.38 103.08 57.38 101.72 58.08 101.72 58.08 103.08 58.76 103.08 58.76 101.72 59.46 101.72 59.46 103.08 59.68 103.08 59.68 101.72 60.38 101.72 60.38 103.08 60.6 103.08 60.6 101.72 61.3 101.72 61.3 103.08 61.98 103.08 61.98 101.72 62.68 101.72 62.68 103.08 63.36 103.08 63.36 101.72 64.06 101.72 64.06 103.08 64.28 103.08 64.28 101.72 64.98 101.72 64.98 103.08 65.66 103.08 65.66 101.72 66.36 101.72 66.36 103.08 67.04 103.08 67.04 101.72 67.74 101.72 67.74 103.08 68.42 103.08 68.42 101.72 69.12 101.72 69.12 103.08 69.34 103.08 69.34 101.72 70.96 101.72 70.96 103.08 72.56 103.08 72.56 101.72 75.56 101.72 75.56 103.08 75.78 103.08 75.78 101.72 76.48 101.72 76.48 103.08 77.16 103.08 77.16 101.72 77.86 101.72 77.86 103.08 78.54 103.08 78.54 101.72 79.24 101.72 79.24 103.08 80.38 103.08 80.38 101.72 81.08 101.72 81.08 103.08 81.76 103.08 81.76 101.72 82.46 101.72 82.46 103.08 83.14 103.08 83.14 101.72 83.84 101.72 83.84 103.08 84.52 103.08 84.52 101.72 85.22 101.72 85.22 103.08 85.9 103.08 85.9 101.72 86.6 101.72 86.6 103.08 87.28 103.08 87.28 101.72 87.98 101.72 87.98 103.08 89.12 103.08 89.12 101.72 89.82 101.72 89.82 103.08 90.5 103.08 90.5 101.72 91.2 101.72 91.2 103.08 91.88 103.08 91.88 101.72 92.58 101.72 92.58 103.08 94.18 103.08 94.18 101.72 94.88 101.72 94.88 103.08 95.56 103.08 95.56 101.72 96.26 101.72 96.26 103.08 96.94 103.08 96.94 101.72 97.64 101.72 97.64 103.08 98.32 103.08 98.32 101.72 99.02 101.72 99.02 103.08 99.7 103.08 99.7 101.72 100.4 101.72 100.4 103.08 101.08 103.08 101.08 101.72 101.78 101.72 101.78 103.08 104.3 103.08 104.3 101.72 105 101.72 105 103.08 105.68 103.08 105.68 101.72 106.38 101.72 106.38 103.08 ;
    LAYER met4 ;
      RECT 139.01 78.29 140.19 79.47 ;
      RECT -0.35 78.29 0.83 79.47 ;
      RECT 139.01 53.99 140.19 55.17 ;
      RECT -0.35 53.99 0.83 55.17 ;
      RECT 139.01 34.77 140.19 35.95 ;
      RECT -0.35 34.77 0.83 35.95 ;
      RECT 139.01 10.29 140.19 11.47 ;
      RECT -0.35 10.29 0.83 11.47 ;
      POLYGON 108.16 102.96 108.16 86.64 125.81 86.64 125.81 85.14 128.11 85.14 128.11 86.64 139.44 86.64 139.44 0.4 128.11 0.4 128.11 1.9 125.81 1.9 125.81 0.4 104.11 0.4 104.11 1.9 101.81 1.9 101.81 0.4 88.49 0.4 88.49 1.9 86.19 1.9 86.19 0.4 76.45 0.4 76.45 1.76 75.35 1.76 75.35 0.4 72.87 0.4 72.87 1.9 70.57 1.9 70.57 0.4 70.01 0.4 70.01 1.2 68.91 1.2 68.91 0.4 57.25 0.4 57.25 1.9 54.95 1.9 54.95 0.4 41.63 0.4 41.63 1.9 39.33 1.9 39.33 0.4 21.23 0.4 21.23 1.9 18.93 1.9 18.93 0.4 5.61 0.4 5.61 1.9 3.31 1.9 3.31 0.4 0.4 0.4 0.4 86.64 3.31 86.64 3.31 85.14 5.61 85.14 5.61 86.64 18.93 86.64 18.93 85.14 21.23 85.14 21.23 86.64 31.68 86.64 31.68 102.96 36.71 102.96 36.71 101.6 37.81 101.6 37.81 102.96 39.33 102.96 39.33 101.46 41.63 101.46 41.63 102.96 44.99 102.96 44.99 101.6 46.09 101.6 46.09 102.96 47.75 102.96 47.75 101.6 48.85 101.6 48.85 102.96 51.43 102.96 51.43 101.6 52.53 101.6 52.53 102.96 54.95 102.96 54.95 101.46 57.25 101.46 57.25 102.96 58.79 102.96 58.79 101.6 59.89 101.6 59.89 102.96 61.55 102.96 61.55 101.6 62.65 101.6 62.65 102.96 65.23 102.96 65.23 101.6 66.33 101.6 66.33 102.96 68.91 102.96 68.91 102.16 70.01 102.16 70.01 102.96 70.57 102.96 70.57 101.46 72.87 101.46 72.87 102.96 74.43 102.96 74.43 101.6 75.53 101.6 75.53 102.96 78.11 102.96 78.11 101.6 79.21 101.6 79.21 102.96 80.87 102.96 80.87 101.6 81.97 101.6 81.97 102.96 83.63 102.96 83.63 101.6 84.73 101.6 84.73 102.96 86.19 102.96 86.19 101.46 88.49 101.46 88.49 102.96 90.07 102.96 90.07 101.6 91.17 101.6 91.17 102.96 92.83 102.96 92.83 101.6 93.93 101.6 93.93 102.96 95.59 102.96 95.59 101.6 96.69 101.6 96.69 102.96 98.35 102.96 98.35 101.6 99.45 101.6 99.45 102.96 101.81 102.96 101.81 101.46 104.11 101.46 104.11 102.96 ;
    LAYER met3 ;
      POLYGON 103.525 103.405 103.525 103.4 103.55 103.4 103.55 103.08 103.525 103.08 103.525 103.075 102.395 103.075 102.395 103.08 102.37 103.08 102.37 103.4 102.395 103.4 102.395 103.405 ;
      POLYGON 72.285 103.405 72.285 103.4 72.31 103.4 72.31 103.08 72.285 103.08 72.285 103.075 71.155 103.075 71.155 103.08 71.13 103.08 71.13 103.4 71.155 103.4 71.155 103.405 ;
      POLYGON 41.045 103.405 41.045 103.4 41.07 103.4 41.07 103.08 41.045 103.08 41.045 103.075 39.915 103.075 39.915 103.08 39.89 103.08 39.89 103.4 39.915 103.4 39.915 103.405 ;
      POLYGON 127.525 87.085 127.525 87.08 127.55 87.08 127.55 86.76 127.525 86.76 127.525 86.755 126.395 86.755 126.395 86.76 126.37 86.76 126.37 87.08 126.395 87.08 126.395 87.085 ;
      POLYGON 20.645 87.085 20.645 87.08 20.67 87.08 20.67 86.76 20.645 86.76 20.645 86.755 19.515 86.755 19.515 86.76 19.49 86.76 19.49 87.08 19.515 87.08 19.515 87.085 ;
      POLYGON 139.765 79.045 139.765 79.04 139.98 79.04 139.98 78.72 139.765 78.72 139.765 78.715 139.435 78.715 139.435 78.72 139.22 78.72 139.22 79.04 139.435 79.04 139.435 79.045 ;
      POLYGON 0.405 79.045 0.405 79.04 0.62 79.04 0.62 78.72 0.405 78.72 0.405 78.715 0.075 78.715 0.075 78.72 -0.14 78.72 -0.14 79.04 0.075 79.04 0.075 79.045 ;
      POLYGON 139.765 54.745 139.765 54.74 139.98 54.74 139.98 54.42 139.765 54.42 139.765 54.415 139.435 54.415 139.435 54.42 139.22 54.42 139.22 54.74 139.435 54.74 139.435 54.745 ;
      POLYGON 0.405 54.745 0.405 54.74 0.62 54.74 0.62 54.42 0.405 54.42 0.405 54.415 0.075 54.415 0.075 54.42 -0.14 54.42 -0.14 54.74 0.075 54.74 0.075 54.745 ;
      POLYGON 139.765 35.525 139.765 35.52 139.98 35.52 139.98 35.2 139.765 35.2 139.765 35.195 139.435 35.195 139.435 35.2 139.22 35.2 139.22 35.52 139.435 35.52 139.435 35.525 ;
      POLYGON 0.405 35.525 0.405 35.52 0.62 35.52 0.62 35.2 0.405 35.2 0.405 35.195 0.075 35.195 0.075 35.2 -0.14 35.2 -0.14 35.52 0.075 35.52 0.075 35.525 ;
      POLYGON 139.765 11.045 139.765 11.04 139.98 11.04 139.98 10.72 139.765 10.72 139.765 10.715 139.435 10.715 139.435 10.72 139.22 10.72 139.22 11.04 139.435 11.04 139.435 11.045 ;
      POLYGON 0.405 11.045 0.405 11.04 0.62 11.04 0.62 10.72 0.405 10.72 0.405 10.715 0.075 10.715 0.075 10.72 -0.14 10.72 -0.14 11.04 0.075 11.04 0.075 11.045 ;
      POLYGON 127.525 0.285 127.525 0.28 127.55 0.28 127.55 -0.04 127.525 -0.04 127.525 -0.045 126.395 -0.045 126.395 -0.04 126.37 -0.04 126.37 0.28 126.395 0.28 126.395 0.285 ;
      POLYGON 103.525 0.285 103.525 0.28 103.55 0.28 103.55 -0.04 103.525 -0.04 103.525 -0.045 102.395 -0.045 102.395 -0.04 102.37 -0.04 102.37 0.28 102.395 0.28 102.395 0.285 ;
      POLYGON 72.285 0.285 72.285 0.28 72.31 0.28 72.31 -0.04 72.285 -0.04 72.285 -0.045 71.155 -0.045 71.155 -0.04 71.13 -0.04 71.13 0.28 71.155 0.28 71.155 0.285 ;
      POLYGON 41.045 0.285 41.045 0.28 41.07 0.28 41.07 -0.04 41.045 -0.04 41.045 -0.045 39.915 -0.045 39.915 -0.04 39.89 -0.04 39.89 0.28 39.915 0.28 39.915 0.285 ;
      POLYGON 20.645 0.285 20.645 0.28 20.67 0.28 20.67 -0.04 20.645 -0.04 20.645 -0.045 19.515 -0.045 19.515 -0.04 19.49 -0.04 19.49 0.28 19.515 0.28 19.515 0.285 ;
      POLYGON 108.16 102.96 108.16 86.64 139.44 86.64 139.44 83.17 138.06 83.17 138.06 82.07 139.44 82.07 139.44 81.13 138.06 81.13 138.06 80.03 139.44 80.03 139.44 77.73 138.06 77.73 138.06 76.63 139.44 76.63 139.44 75.69 138.06 75.69 138.06 74.59 139.44 74.59 139.44 73.65 138.06 73.65 138.06 72.55 139.44 72.55 139.44 71.61 138.06 71.61 138.06 70.51 139.44 70.51 139.44 69.57 138.06 69.57 138.06 68.47 139.44 68.47 139.44 67.53 138.06 67.53 138.06 66.43 139.44 66.43 139.44 65.49 138.06 65.49 138.06 64.39 139.44 64.39 139.44 62.09 138.06 62.09 138.06 60.99 139.44 60.99 139.44 59.37 138.06 59.37 138.06 58.27 139.44 58.27 139.44 57.33 138.06 57.33 138.06 56.23 139.44 56.23 139.44 53.25 138.06 53.25 138.06 52.15 139.44 52.15 139.44 51.21 138.06 51.21 138.06 50.11 139.44 50.11 139.44 49.17 138.06 49.17 138.06 48.07 139.44 48.07 139.44 47.13 138.06 47.13 138.06 46.03 139.44 46.03 139.44 45.09 138.06 45.09 138.06 43.99 139.44 43.99 139.44 43.05 138.06 43.05 138.06 41.95 139.44 41.95 139.44 41.01 138.06 41.01 138.06 39.91 139.44 39.91 139.44 38.97 138.06 38.97 138.06 37.87 139.44 37.87 139.44 36.93 138.06 36.93 138.06 35.83 139.44 35.83 139.44 34.21 138.06 34.21 138.06 33.11 139.44 33.11 139.44 32.17 138.06 32.17 138.06 31.07 139.44 31.07 139.44 30.13 138.06 30.13 138.06 29.03 139.44 29.03 139.44 28.09 138.06 28.09 138.06 26.99 139.44 26.99 139.44 21.97 138.06 21.97 138.06 20.87 139.44 20.87 139.44 19.93 138.06 19.93 138.06 18.83 139.44 18.83 139.44 17.89 138.06 17.89 138.06 16.79 139.44 16.79 139.44 15.85 138.06 15.85 138.06 14.75 139.44 14.75 139.44 13.81 138.06 13.81 138.06 12.71 139.44 12.71 139.44 9.73 138.06 9.73 138.06 8.63 139.44 8.63 139.44 7.69 138.06 7.69 138.06 6.59 139.44 6.59 139.44 5.65 138.06 5.65 138.06 4.55 139.44 4.55 139.44 4.29 138.06 4.29 138.06 3.19 139.44 3.19 139.44 0.4 0.4 0.4 0.4 3.87 1.78 3.87 1.78 4.97 0.4 4.97 0.4 5.23 1.78 5.23 1.78 6.33 0.4 6.33 0.4 6.59 1.78 6.59 1.78 7.69 0.4 7.69 0.4 7.95 1.78 7.95 1.78 9.05 0.4 9.05 0.4 9.31 1.78 9.31 1.78 10.41 0.4 10.41 0.4 12.71 1.78 12.71 1.78 13.81 0.4 13.81 0.4 14.75 1.78 14.75 1.78 15.85 0.4 15.85 0.4 16.79 1.78 16.79 1.78 17.89 0.4 17.89 0.4 18.83 1.78 18.83 1.78 19.93 0.4 19.93 0.4 20.87 1.78 20.87 1.78 21.97 0.4 21.97 0.4 22.91 1.78 22.91 1.78 24.01 0.4 24.01 0.4 24.95 1.78 24.95 1.78 26.05 0.4 26.05 0.4 26.99 1.78 26.99 1.78 28.09 0.4 28.09 0.4 29.03 1.78 29.03 1.78 30.13 0.4 30.13 0.4 31.07 1.78 31.07 1.78 32.17 0.4 32.17 0.4 33.11 1.78 33.11 1.78 34.21 0.4 34.21 0.4 35.83 1.78 35.83 1.78 36.93 0.4 36.93 0.4 37.87 1.78 37.87 1.78 38.97 0.4 38.97 0.4 39.91 1.78 39.91 1.78 41.01 0.4 41.01 0.4 41.95 1.78 41.95 1.78 43.05 0.4 43.05 0.4 43.99 1.78 43.99 1.78 45.09 0.4 45.09 0.4 46.03 1.78 46.03 1.78 47.13 0.4 47.13 0.4 48.07 1.78 48.07 1.78 49.17 0.4 49.17 0.4 50.11 1.78 50.11 1.78 51.21 0.4 51.21 0.4 52.15 1.78 52.15 1.78 53.25 0.4 53.25 0.4 56.23 1.78 56.23 1.78 57.33 0.4 57.33 0.4 58.27 1.78 58.27 1.78 59.37 0.4 59.37 0.4 60.31 1.78 60.31 1.78 61.41 0.4 61.41 0.4 62.35 1.78 62.35 1.78 63.45 0.4 63.45 0.4 64.39 1.78 64.39 1.78 65.49 0.4 65.49 0.4 67.11 1.78 67.11 1.78 68.21 0.4 68.21 0.4 69.15 1.78 69.15 1.78 70.25 0.4 70.25 0.4 71.19 1.78 71.19 1.78 72.29 0.4 72.29 0.4 73.23 1.78 73.23 1.78 74.33 0.4 74.33 0.4 75.27 1.78 75.27 1.78 76.37 0.4 76.37 0.4 77.31 1.78 77.31 1.78 78.41 0.4 78.41 0.4 80.03 1.78 80.03 1.78 81.13 0.4 81.13 0.4 82.07 1.78 82.07 1.78 83.17 0.4 83.17 0.4 86.64 31.68 86.64 31.68 95.67 33.06 95.67 33.06 96.77 31.68 96.77 31.68 102.96 ;
    LAYER met1 ;
      POLYGON 107.8 103.6 107.8 103.12 103.6 103.12 103.6 103.11 102.32 103.11 102.32 103.12 72.36 103.12 72.36 103.11 71.08 103.11 71.08 103.12 41.12 103.12 41.12 103.11 39.84 103.11 39.84 103.12 32.04 103.12 32.04 103.6 ;
      POLYGON 139.08 87.28 139.08 86.8 127.6 86.8 127.6 86.79 126.32 86.79 126.32 86.8 20.72 86.8 20.72 86.79 19.44 86.79 19.44 86.8 0.76 86.8 0.76 87.28 ;
      POLYGON 127.6 0.25 127.6 0.24 139.08 0.24 139.08 -0.24 0.76 -0.24 0.76 0.24 19.44 0.24 19.44 0.25 20.72 0.25 20.72 0.24 39.84 0.24 39.84 0.25 41.12 0.25 41.12 0.24 71.08 0.24 71.08 0.25 72.36 0.25 72.36 0.24 102.32 0.24 102.32 0.25 103.6 0.25 103.6 0.24 126.32 0.24 126.32 0.25 ;
      POLYGON 107.8 103.08 107.8 102.84 108.28 102.84 108.28 101.16 107.8 101.16 107.8 100.12 108.28 100.12 108.28 98.44 107.8 98.44 107.8 97.4 108.28 97.4 108.28 95.72 107.8 95.72 107.8 94.68 108.28 94.68 108.28 93 107.8 93 107.8 91.96 108.28 91.96 108.28 90.28 107.8 90.28 107.8 89.24 108.28 89.24 108.28 86.76 139.08 86.76 139.08 86.52 139.56 86.52 139.56 85.52 138.965 85.52 138.965 84.82 139.08 84.82 139.08 83.8 139.56 83.8 139.56 83.14 138.965 83.14 138.965 82.44 139.56 82.44 139.56 82.12 139.08 82.12 139.08 81.1 138.965 81.1 138.965 79.72 139.56 79.72 139.56 79.4 139.08 79.4 139.08 78.38 138.965 78.38 138.965 77 139.56 77 139.56 76.68 139.08 76.68 139.08 75.66 138.965 75.66 138.965 74.28 139.56 74.28 139.56 73.96 139.08 73.96 139.08 72.92 139.56 72.92 139.56 72.26 138.965 72.26 138.965 71.56 139.56 71.56 139.56 71.24 139.08 71.24 139.08 70.2 139.56 70.2 139.56 69.54 138.965 69.54 138.965 68.84 139.56 68.84 139.56 68.52 139.08 68.52 139.08 67.48 139.56 67.48 139.56 66.82 138.965 66.82 138.965 66.12 139.56 66.12 139.56 65.8 139.08 65.8 139.08 64.76 139.56 64.76 139.56 64.44 138.965 64.44 138.965 63.74 139.56 63.74 139.56 63.08 139.08 63.08 139.08 62.04 139.56 62.04 139.56 61.38 138.965 61.38 138.965 60.68 139.56 60.68 139.56 60.36 139.08 60.36 139.08 59.32 139.56 59.32 139.56 58.66 138.965 58.66 138.965 57.96 139.56 57.96 139.56 57.64 139.08 57.64 139.08 56.6 139.56 56.6 139.56 56.28 138.965 56.28 138.965 55.58 139.56 55.58 139.56 54.92 139.08 54.92 139.08 53.88 139.56 53.88 139.56 53.56 138.965 53.56 138.965 52.86 139.56 52.86 139.56 52.2 139.08 52.2 139.08 51.16 139.56 51.16 139.56 50.84 138.965 50.84 138.965 50.14 139.56 50.14 139.56 49.48 139.08 49.48 139.08 48.44 139.56 48.44 139.56 48.12 138.965 48.12 138.965 47.42 139.56 47.42 139.56 46.76 139.08 46.76 139.08 45.72 139.56 45.72 139.56 45.06 138.965 45.06 138.965 44.36 139.56 44.36 139.56 44.04 139.08 44.04 139.08 43 139.56 43 139.56 42.34 138.965 42.34 138.965 41.64 139.56 41.64 139.56 41.32 139.08 41.32 139.08 40.28 139.56 40.28 139.56 39.62 138.965 39.62 138.965 38.92 139.56 38.92 139.56 38.6 139.08 38.6 139.08 37.56 139.56 37.56 139.56 37.24 138.965 37.24 138.965 35.86 139.08 35.86 139.08 34.84 139.56 34.84 139.56 34.52 138.965 34.52 138.965 33.14 139.08 33.14 139.08 32.12 139.56 32.12 139.56 31.46 138.965 31.46 138.965 30.76 139.56 30.76 139.56 30.44 139.08 30.44 139.08 29.4 139.56 29.4 139.56 29.08 138.965 29.08 138.965 28.38 139.56 28.38 139.56 27.72 139.08 27.72 139.08 26.68 139.56 26.68 139.56 26.36 138.965 26.36 138.965 25.66 139.56 25.66 139.56 25 139.08 25 139.08 23.96 139.56 23.96 139.56 23.64 138.965 23.64 138.965 22.94 139.56 22.94 139.56 22.28 139.08 22.28 139.08 21.24 139.56 21.24 139.56 20.92 138.965 20.92 138.965 20.22 139.56 20.22 139.56 19.56 139.08 19.56 139.08 18.52 139.56 18.52 139.56 17.86 138.965 17.86 138.965 17.16 139.56 17.16 139.56 16.84 139.08 16.84 139.08 15.8 139.56 15.8 139.56 15.48 138.965 15.48 138.965 14.1 139.08 14.1 139.08 13.08 139.56 13.08 139.56 12.76 138.965 12.76 138.965 12.06 139.56 12.06 139.56 11.4 139.08 11.4 139.08 10.36 139.56 10.36 139.56 10.04 138.965 10.04 138.965 9.34 139.56 9.34 139.56 8.68 139.08 8.68 139.08 7.64 139.56 7.64 139.56 7.32 138.965 7.32 138.965 6.62 139.56 6.62 139.56 5.96 139.08 5.96 139.08 4.92 139.56 4.92 139.56 4.6 138.965 4.6 138.965 3.9 139.56 3.9 139.56 3.24 139.08 3.24 139.08 2.22 138.965 2.22 138.965 1.52 139.56 1.52 139.56 0.52 139.08 0.52 139.08 0.28 0.76 0.28 0.76 0.52 0.28 0.52 0.28 1.52 0.875 1.52 0.875 2.22 0.76 2.22 0.76 3.24 0.28 3.24 0.28 3.9 0.875 3.9 0.875 4.6 0.28 4.6 0.28 4.92 0.76 4.92 0.76 5.96 0.28 5.96 0.28 6.62 0.875 6.62 0.875 7.32 0.28 7.32 0.28 7.64 0.76 7.64 0.76 8.68 0.28 8.68 0.28 9.34 0.875 9.34 0.875 10.04 0.28 10.04 0.28 10.36 0.76 10.36 0.76 11.4 0.28 11.4 0.28 12.06 0.875 12.06 0.875 12.76 0.28 12.76 0.28 13.08 0.76 13.08 0.76 14.12 0.28 14.12 0.28 14.78 0.875 14.78 0.875 15.48 0.28 15.48 0.28 15.8 0.76 15.8 0.76 16.84 0.28 16.84 0.28 17.16 0.875 17.16 0.875 18.54 0.76 18.54 0.76 19.56 0.28 19.56 0.28 20.22 0.875 20.22 0.875 20.92 0.28 20.92 0.28 21.24 0.76 21.24 0.76 22.28 0.28 22.28 0.28 22.94 0.875 22.94 0.875 23.64 0.28 23.64 0.28 23.96 0.76 23.96 0.76 25 0.28 25 0.28 25.66 0.875 25.66 0.875 26.36 0.28 26.36 0.28 26.68 0.76 26.68 0.76 27.72 0.28 27.72 0.28 28.38 0.875 28.38 0.875 29.08 0.28 29.08 0.28 29.4 0.76 29.4 0.76 30.44 0.28 30.44 0.28 31.1 0.875 31.1 0.875 31.8 0.28 31.8 0.28 32.12 0.76 32.12 0.76 33.16 0.28 33.16 0.28 33.82 0.875 33.82 0.875 34.52 0.28 34.52 0.28 34.84 0.76 34.84 0.76 35.86 0.875 35.86 0.875 37.24 0.28 37.24 0.28 37.56 0.76 37.56 0.76 38.6 0.28 38.6 0.28 38.92 0.875 38.92 0.875 39.62 0.28 39.62 0.28 40.28 0.76 40.28 0.76 41.32 0.28 41.32 0.28 41.64 0.875 41.64 0.875 42.34 0.28 42.34 0.28 43 0.76 43 0.76 44.04 0.28 44.04 0.28 44.36 0.875 44.36 0.875 45.06 0.28 45.06 0.28 45.72 0.76 45.72 0.76 46.76 0.28 46.76 0.28 47.42 0.875 47.42 0.875 48.12 0.28 48.12 0.28 48.44 0.76 48.44 0.76 49.48 0.28 49.48 0.28 50.14 0.875 50.14 0.875 50.84 0.28 50.84 0.28 51.16 0.76 51.16 0.76 52.2 0.28 52.2 0.28 52.52 0.875 52.52 0.875 53.22 0.28 53.22 0.28 53.88 0.76 53.88 0.76 54.9 0.875 54.9 0.875 56.28 0.28 56.28 0.28 56.6 0.76 56.6 0.76 57.64 0.28 57.64 0.28 57.96 0.875 57.96 0.875 58.66 0.28 58.66 0.28 59.32 0.76 59.32 0.76 60.36 0.28 60.36 0.28 60.68 0.875 60.68 0.875 61.38 0.28 61.38 0.28 62.04 0.76 62.04 0.76 63.08 0.28 63.08 0.28 63.4 0.875 63.4 0.875 64.1 0.28 64.1 0.28 64.76 0.76 64.76 0.76 65.8 0.28 65.8 0.28 66.12 0.875 66.12 0.875 66.82 0.28 66.82 0.28 67.48 0.76 67.48 0.76 68.52 0.28 68.52 0.28 68.84 0.875 68.84 0.875 69.54 0.28 69.54 0.28 70.2 0.76 70.2 0.76 71.24 0.28 71.24 0.28 71.56 0.875 71.56 0.875 72.26 0.28 72.26 0.28 72.92 0.76 72.92 0.76 73.96 0.28 73.96 0.28 74.28 0.875 74.28 0.875 74.98 0.28 74.98 0.28 75.64 0.76 75.64 0.76 76.68 0.28 76.68 0.28 77 0.875 77 0.875 77.7 0.28 77.7 0.28 78.36 0.76 78.36 0.76 79.4 0.28 79.4 0.28 79.72 0.875 79.72 0.875 80.42 0.28 80.42 0.28 81.08 0.76 81.08 0.76 82.12 0.28 82.12 0.28 82.44 0.875 82.44 0.875 83.14 0.28 83.14 0.28 83.8 0.76 83.8 0.76 84.84 0.28 84.84 0.28 86.52 0.76 86.52 0.76 86.76 31.56 86.76 31.56 89.24 32.04 89.24 32.04 90.28 31.56 90.28 31.56 91.96 32.04 91.96 32.04 93 31.56 93 31.56 94.68 32.04 94.68 32.04 95.72 31.56 95.72 31.56 96.04 32.155 96.04 32.155 97.42 32.04 97.42 32.04 98.44 31.56 98.44 31.56 100.12 32.04 100.12 32.04 101.16 31.56 101.16 31.56 102.84 32.04 102.84 32.04 103.08 ;
    LAYER met5 ;
      RECT 138.8 52.18 140.4 52.92 ;
      RECT -0.56 52.18 1.04 52.92 ;
      RECT 138.8 8.48 140.4 8.92 ;
      RECT -0.56 8.48 1.04 8.92 ;
      POLYGON 106.96 101.76 106.96 85.44 138.24 85.44 138.24 82.92 133.44 82.92 133.44 74.92 138.24 74.92 138.24 60.92 133.44 60.92 133.44 52.92 138.24 52.92 138.24 38.92 133.44 38.92 133.44 30.92 138.24 30.92 138.24 16.92 133.44 16.92 133.44 8.92 138.24 8.92 138.24 1.6 1.6 1.6 1.6 8.92 6.4 8.92 6.4 16.92 1.6 16.92 1.6 30.92 6.4 30.92 6.4 38.92 1.6 38.92 1.6 52.92 6.4 52.92 6.4 60.92 1.6 60.92 1.6 74.92 6.4 74.92 6.4 82.92 1.6 82.92 1.6 85.44 32.88 85.44 32.88 101.76 ;
    LAYER li1 ;
      POLYGON 108.56 103.445 108.56 103.275 108.015 103.275 108.015 101.665 106.805 101.665 106.805 102.185 105.425 102.185 105.425 103.275 104.745 103.275 104.745 102.135 104.575 102.135 104.575 103.275 102.205 103.275 102.205 102.515 102.035 102.515 102.035 103.275 100.655 103.275 100.655 101.665 99.905 101.665 99.905 102.185 98.985 102.185 98.985 103.275 98.815 103.275 98.815 102.11 98.525 102.11 98.525 103.275 97.925 103.275 97.925 102.135 97.62 102.135 97.62 103.275 97.28 103.275 97.28 102.895 96.95 102.895 96.95 103.275 96.43 103.275 96.43 102.815 96.18 102.815 96.18 103.275 94.565 103.275 94.565 102.815 94.195 102.815 94.195 103.275 93.56 103.275 93.56 102.845 93.23 102.845 93.23 103.275 91.34 103.275 91.34 102.815 91.09 102.815 91.09 103.275 90.085 103.275 90.085 102.775 89.755 102.775 89.755 103.275 89.155 103.275 89.155 101.645 88.635 101.645 88.635 102.185 87.945 102.185 87.945 103.275 87.775 103.275 87.775 101.665 86.085 101.665 86.085 102.185 84.265 102.185 84.265 103.275 84.095 103.275 84.095 102.11 83.805 102.11 83.805 103.275 83.125 103.275 83.125 102.135 82.955 102.135 82.955 103.275 80.585 103.275 80.585 102.515 80.415 102.515 80.415 103.275 79.495 103.275 79.495 101.665 78.745 101.665 78.745 102.185 77.825 102.185 77.825 103.275 76.905 103.275 76.905 102.515 76.735 102.515 76.735 103.275 74.365 103.275 74.365 102.135 74.195 102.135 74.195 103.275 73.055 103.275 73.055 101.665 71.365 101.665 71.365 102.185 69.545 102.185 69.545 103.275 69.375 103.275 69.375 102.11 69.085 102.11 69.085 103.275 68.455 103.275 68.455 101.665 67.245 101.665 67.245 102.185 65.865 102.185 65.865 103.275 65.69 103.275 65.69 101.665 63.095 101.665 63.095 102.185 60.345 102.185 60.345 103.275 60.17 103.275 60.17 101.665 57.575 101.665 57.575 102.185 54.825 102.185 54.825 103.275 54.655 103.275 54.655 102.11 54.365 102.11 54.365 103.275 53.685 103.275 53.685 102.135 53.515 102.135 53.515 103.275 51.145 103.275 51.145 102.515 50.975 102.515 50.975 103.275 49.595 103.275 49.595 101.665 48.845 101.665 48.845 102.185 47.925 102.185 47.925 103.275 47.245 103.275 47.245 102.135 47.075 102.135 47.075 103.275 44.705 103.275 44.705 102.515 44.535 102.515 44.535 103.275 43.615 103.275 43.615 101.665 41.925 101.665 41.925 102.185 40.105 102.185 40.105 103.275 39.935 103.275 39.935 102.11 39.645 102.11 39.645 103.275 38.965 103.275 38.965 102.135 38.795 102.135 38.795 103.275 36.425 103.275 36.425 102.515 36.255 102.515 36.255 103.275 34.875 103.275 34.875 101.665 33.185 101.665 33.185 102.185 31.365 102.185 31.365 103.275 31.28 103.275 31.28 103.445 ;
      POLYGON 33.015 102.015 33.015 101.495 34.875 101.495 34.875 100.725 36.8 100.725 36.8 100.555 36.71 100.555 36.71 99.785 33.945 99.785 33.945 99.265 31.365 99.265 31.365 100.555 31.28 100.555 31.28 100.725 31.365 100.725 31.365 102.015 ;
      RECT 108.1 100.555 108.56 100.725 ;
      POLYGON 36.71 99.615 36.71 98.005 36.8 98.005 36.8 97.835 34.875 97.835 34.875 96.225 33.185 96.225 33.185 96.745 31.365 96.745 31.365 97.835 31.28 97.835 31.28 98.005 31.365 98.005 31.365 99.095 34.115 99.095 34.115 99.615 ;
      RECT 108.1 97.835 108.56 98.005 ;
      POLYGON 33.015 96.575 33.015 96.055 34.875 96.055 34.875 95.285 36.8 95.285 36.8 95.115 36.71 95.115 36.71 94.345 33.945 94.345 33.945 93.825 31.365 93.825 31.365 95.115 31.28 95.115 31.28 95.285 31.365 95.285 31.365 96.575 ;
      RECT 108.1 95.115 108.56 95.285 ;
      POLYGON 36.71 94.175 36.71 92.565 36.8 92.565 36.8 92.395 33.955 92.395 33.955 90.785 32.745 90.785 32.745 91.305 31.365 91.305 31.365 92.395 31.28 92.395 31.28 92.565 31.365 92.565 31.365 93.655 34.115 93.655 34.115 94.175 ;
      RECT 108.1 92.395 108.56 92.565 ;
      POLYGON 32.575 91.135 32.575 90.615 33.955 90.615 33.955 89.845 34.96 89.845 34.96 89.675 34.875 89.675 34.875 88.905 33.015 88.905 33.015 88.385 31.365 88.385 31.365 89.675 31.28 89.675 31.28 89.845 31.365 89.845 31.365 91.135 ;
      RECT 108.1 89.675 108.56 89.845 ;
      POLYGON 34.875 88.735 34.875 87.125 34.96 87.125 34.96 86.955 33.985 86.955 33.985 85.815 33.68 85.815 33.68 86.955 33.34 86.955 33.34 86.575 33.01 86.575 33.01 86.955 32.49 86.955 32.49 86.495 32.24 86.495 32.24 86.955 30.625 86.955 30.625 86.495 30.255 86.495 30.255 86.955 29.62 86.955 29.62 86.525 29.29 86.525 29.29 86.955 27.4 86.955 27.4 86.495 27.15 86.495 27.15 86.955 26.145 86.955 26.145 86.455 25.815 86.455 25.815 86.955 25.215 86.955 25.215 85.79 24.925 85.79 24.925 86.955 24.755 86.955 24.755 85.325 24.235 85.325 24.235 85.865 23.545 85.865 23.545 86.955 23.375 86.955 23.375 85.345 21.685 85.345 21.685 85.865 19.865 85.865 19.865 86.955 19.265 86.955 19.265 85.815 18.96 85.815 18.96 86.955 18.62 86.955 18.62 86.575 18.29 86.575 18.29 86.955 17.77 86.955 17.77 86.495 17.52 86.495 17.52 86.955 15.905 86.955 15.905 86.495 15.535 86.495 15.535 86.955 14.9 86.955 14.9 86.525 14.57 86.525 14.57 86.955 12.68 86.955 12.68 86.495 12.43 86.495 12.43 86.955 11.425 86.955 11.425 86.455 11.095 86.455 11.095 86.955 10.495 86.955 10.495 85.79 10.205 85.79 10.205 86.955 9.115 86.955 9.115 85.345 7.425 85.345 7.425 85.865 5.605 85.865 5.605 86.955 5.43 86.955 5.43 85.345 2.835 85.345 2.835 85.865 0.085 85.865 0.085 86.955 0 86.955 0 87.125 31.365 87.125 31.365 88.215 33.185 88.215 33.185 88.735 ;
      POLYGON 139.84 87.125 139.84 86.955 139.295 86.955 139.295 85.345 137.605 85.345 137.605 85.865 135.785 85.865 135.785 86.955 135.615 86.955 135.615 85.79 135.325 85.79 135.325 86.955 135.155 86.955 135.155 85.345 133.945 85.345 133.945 85.865 132.565 85.865 132.565 86.955 131.885 86.955 131.885 85.815 131.715 85.815 131.715 86.955 129.345 86.955 129.345 86.195 129.175 86.195 129.175 86.955 128.255 86.955 128.255 85.79 127.965 85.79 127.965 86.955 127.335 86.955 127.335 85.345 125.645 85.345 125.645 85.865 123.825 85.865 123.825 86.955 123.145 86.955 123.145 86.155 122.975 86.155 122.975 86.955 122.305 86.955 122.305 86.155 122.135 86.155 122.135 86.955 121.545 86.955 121.545 86.155 121.215 86.155 121.215 86.955 120.705 86.955 120.705 86.155 120.375 86.155 120.375 86.955 119.865 86.955 119.865 86.155 119.535 86.155 119.535 86.955 119.025 86.955 119.025 85.805 118.695 85.805 118.695 86.955 117.215 86.955 117.215 85.345 115.525 85.345 115.525 85.865 113.705 85.865 113.705 86.955 113.535 86.955 113.535 85.79 113.245 85.79 113.245 86.955 112.645 86.955 112.645 85.815 112.34 85.815 112.34 86.955 112 86.955 112 86.575 111.67 86.575 111.67 86.955 111.15 86.955 111.15 86.495 110.9 86.495 110.9 86.955 109.285 86.955 109.285 86.495 108.915 86.495 108.915 86.955 108.28 86.955 108.28 86.525 107.95 86.525 107.95 86.955 106.06 86.955 106.06 86.495 105.81 86.495 105.81 86.955 104.805 86.955 104.805 86.455 104.475 86.455 104.475 86.955 103.96 86.955 103.96 87.125 ;
      POLYGON 2.665 85.695 2.665 85.175 5.43 85.175 5.43 84.405 5.52 84.405 5.52 84.235 5.43 84.235 5.43 83.465 2.665 83.465 2.665 82.945 0.085 82.945 0.085 84.235 0 84.235 0 84.405 0.085 84.405 0.085 85.695 ;
      RECT 139.38 84.235 139.84 84.405 ;
      POLYGON 5.43 83.295 5.43 81.685 5.52 81.685 5.52 81.515 2.675 81.515 2.675 79.905 1.465 79.905 1.465 80.425 0.085 80.425 0.085 81.515 0 81.515 0 81.685 0.085 81.685 0.085 82.775 2.835 82.775 2.835 83.295 ;
      RECT 139.38 81.515 139.84 81.685 ;
      POLYGON 1.295 80.255 1.295 79.735 2.675 79.735 2.675 78.965 5.52 78.965 5.52 78.795 5.43 78.795 5.43 78.025 2.665 78.025 2.665 77.505 0.085 77.505 0.085 78.795 0 78.795 0 78.965 0.085 78.965 0.085 80.255 ;
      RECT 139.38 78.795 139.84 78.965 ;
      POLYGON 5.43 77.855 5.43 76.245 5.52 76.245 5.52 76.075 2.675 76.075 2.675 74.465 1.465 74.465 1.465 74.985 0.085 74.985 0.085 76.075 0 76.075 0 76.245 0.085 76.245 0.085 77.335 2.835 77.335 2.835 77.855 ;
      RECT 139.38 76.075 139.84 76.245 ;
      POLYGON 1.295 74.815 1.295 74.295 2.675 74.295 2.675 73.525 5.52 73.525 5.52 73.355 5.43 73.355 5.43 72.585 2.665 72.585 2.665 72.065 0.085 72.065 0.085 73.355 0 73.355 0 73.525 0.085 73.525 0.085 74.815 ;
      RECT 139.38 73.355 139.84 73.525 ;
      POLYGON 5.43 72.415 5.43 70.805 5.52 70.805 5.52 70.635 2.675 70.635 2.675 69.025 1.465 69.025 1.465 69.545 0.085 69.545 0.085 70.635 0 70.635 0 70.805 0.085 70.805 0.085 71.895 2.835 71.895 2.835 72.415 ;
      POLYGON 139.84 70.805 139.84 70.635 139.755 70.635 139.755 69.025 138.545 69.025 138.545 69.545 137.165 69.545 137.165 70.635 137.08 70.635 137.08 70.805 ;
      POLYGON 138.375 69.375 138.375 68.855 139.755 68.855 139.755 68.085 139.84 68.085 139.84 67.915 137.08 67.915 137.08 68.085 137.165 68.085 137.165 69.375 ;
      POLYGON 1.295 69.375 1.295 68.855 2.675 68.855 2.675 68.085 5.52 68.085 5.52 67.915 5.43 67.915 5.43 67.145 2.665 67.145 2.665 66.625 0.085 66.625 0.085 67.915 0 67.915 0 68.085 0.085 68.085 0.085 69.375 ;
      POLYGON 5.43 66.975 5.43 65.365 5.52 65.365 5.52 65.195 3.595 65.195 3.595 63.585 1.905 63.585 1.905 64.105 0.085 64.105 0.085 65.195 0 65.195 0 65.365 0.085 65.365 0.085 66.455 2.835 66.455 2.835 66.975 ;
      POLYGON 139.84 65.365 139.84 65.195 139.755 65.195 139.755 63.585 138.065 63.585 138.065 64.105 136.245 64.105 136.245 65.195 136.16 65.195 136.16 65.365 ;
      POLYGON 137.895 63.935 137.895 63.415 139.755 63.415 139.755 62.645 139.84 62.645 139.84 62.475 136.16 62.475 136.16 62.645 136.245 62.645 136.245 63.935 ;
      POLYGON 1.735 63.935 1.735 63.415 3.595 63.415 3.595 62.645 3.68 62.645 3.68 62.475 3.595 62.475 3.595 61.705 1.735 61.705 1.735 61.185 0.085 61.185 0.085 62.475 0 62.475 0 62.645 0.085 62.645 0.085 63.935 ;
      POLYGON 3.595 61.535 3.595 59.925 5.52 59.925 5.52 59.755 5.43 59.755 5.43 58.145 2.835 58.145 2.835 58.665 0.085 58.665 0.085 59.755 0 59.755 0 59.925 0.085 59.925 0.085 61.015 1.905 61.015 1.905 61.535 ;
      POLYGON 139.84 59.925 139.84 59.755 139.755 59.755 139.755 58.145 138.065 58.145 138.065 58.665 136.245 58.665 136.245 59.755 136.16 59.755 136.16 59.925 ;
      POLYGON 137.895 58.495 137.895 57.975 139.755 57.975 139.755 57.205 139.84 57.205 139.84 57.035 136.16 57.035 136.16 57.205 136.245 57.205 136.245 58.495 ;
      POLYGON 2.665 58.495 2.665 57.975 5.43 57.975 5.43 57.205 5.52 57.205 5.52 57.035 3.595 57.035 3.595 56.265 1.735 56.265 1.735 55.745 0.085 55.745 0.085 57.035 0 57.035 0 57.205 0.085 57.205 0.085 58.495 ;
      POLYGON 3.595 56.095 3.595 54.485 3.68 54.485 3.68 54.315 3.595 54.315 3.595 52.705 1.905 52.705 1.905 53.225 0.085 53.225 0.085 54.315 0 54.315 0 54.485 0.085 54.485 0.085 55.575 1.905 55.575 1.905 56.095 ;
      RECT 139.38 54.315 139.84 54.485 ;
      POLYGON 1.735 53.055 1.735 52.535 3.595 52.535 3.595 51.765 3.68 51.765 3.68 51.595 3.595 51.595 3.595 50.825 1.735 50.825 1.735 50.305 0.085 50.305 0.085 51.595 0 51.595 0 51.765 0.085 51.765 0.085 53.055 ;
      RECT 139.38 51.595 139.84 51.765 ;
      POLYGON 3.595 50.655 3.595 49.045 3.68 49.045 3.68 48.875 3.595 48.875 3.595 47.265 1.905 47.265 1.905 47.785 0.085 47.785 0.085 48.875 0 48.875 0 49.045 0.085 49.045 0.085 50.135 1.905 50.135 1.905 50.655 ;
      RECT 139.38 48.875 139.84 49.045 ;
      POLYGON 1.735 47.615 1.735 47.095 3.595 47.095 3.595 46.325 3.68 46.325 3.68 46.155 3.595 46.155 3.595 45.385 1.735 45.385 1.735 44.865 0.085 44.865 0.085 46.155 0 46.155 0 46.325 0.085 46.325 0.085 47.615 ;
      RECT 139.38 46.155 139.84 46.325 ;
      POLYGON 3.595 45.215 3.595 43.605 5.52 43.605 5.52 43.435 5.43 43.435 5.43 41.825 2.835 41.825 2.835 42.345 0.085 42.345 0.085 43.435 0 43.435 0 43.605 0.085 43.605 0.085 44.695 1.905 44.695 1.905 45.215 ;
      RECT 139.38 43.435 139.84 43.605 ;
      POLYGON 2.665 42.175 2.665 41.655 5.43 41.655 5.43 40.885 5.52 40.885 5.52 40.715 5.43 40.715 5.43 39.945 2.665 39.945 2.665 39.425 0.085 39.425 0.085 40.715 0 40.715 0 40.885 0.085 40.885 0.085 42.175 ;
      RECT 139.38 40.715 139.84 40.885 ;
      POLYGON 5.43 39.775 5.43 38.165 5.52 38.165 5.52 37.995 3.595 37.995 3.595 36.385 1.905 36.385 1.905 36.905 0.085 36.905 0.085 37.995 0 37.995 0 38.165 0.085 38.165 0.085 39.255 2.835 39.255 2.835 39.775 ;
      RECT 139.38 37.995 139.84 38.165 ;
      POLYGON 1.735 36.735 1.735 36.215 3.595 36.215 3.595 35.445 5.52 35.445 5.52 35.275 5.43 35.275 5.43 34.505 2.665 34.505 2.665 33.985 0.085 33.985 0.085 35.275 0 35.275 0 35.445 0.085 35.445 0.085 36.735 ;
      RECT 139.38 35.275 139.84 35.445 ;
      POLYGON 5.43 34.335 5.43 32.725 5.52 32.725 5.52 32.555 5.43 32.555 5.43 30.945 2.835 30.945 2.835 31.465 0.085 31.465 0.085 32.555 0 32.555 0 32.725 0.085 32.725 0.085 33.815 2.835 33.815 2.835 34.335 ;
      RECT 139.38 32.555 139.84 32.725 ;
      POLYGON 2.665 31.295 2.665 30.775 5.43 30.775 5.43 30.005 5.52 30.005 5.52 29.835 5.43 29.835 5.43 29.065 2.665 29.065 2.665 28.545 0.085 28.545 0.085 29.835 0 29.835 0 30.005 0.085 30.005 0.085 31.295 ;
      RECT 139.38 29.835 139.84 30.005 ;
      POLYGON 5.43 28.895 5.43 27.285 5.52 27.285 5.52 27.115 3.595 27.115 3.595 25.505 1.905 25.505 1.905 26.025 0.085 26.025 0.085 27.115 0 27.115 0 27.285 0.085 27.285 0.085 28.375 2.835 28.375 2.835 28.895 ;
      RECT 139.38 27.115 139.84 27.285 ;
      POLYGON 1.735 25.855 1.735 25.335 3.595 25.335 3.595 24.565 5.52 24.565 5.52 24.395 5.43 24.395 5.43 23.625 2.665 23.625 2.665 23.105 0.085 23.105 0.085 24.395 0 24.395 0 24.565 0.085 24.565 0.085 25.855 ;
      RECT 139.38 24.395 139.84 24.565 ;
      POLYGON 5.43 23.455 5.43 21.845 5.52 21.845 5.52 21.675 5.43 21.675 5.43 20.065 2.835 20.065 2.835 20.585 0.085 20.585 0.085 21.675 0 21.675 0 21.845 0.085 21.845 0.085 22.935 2.835 22.935 2.835 23.455 ;
      POLYGON 139.84 21.845 139.84 21.675 139.755 21.675 139.755 20.045 139.235 20.045 139.235 20.585 138.545 20.585 138.545 21.675 138.46 21.675 138.46 21.845 ;
      POLYGON 139.065 20.415 139.065 19.875 139.755 19.875 139.755 19.125 139.84 19.125 139.84 18.955 138.46 18.955 138.46 19.125 138.545 19.125 138.545 20.415 ;
      POLYGON 2.665 20.415 2.665 19.895 5.43 19.895 5.43 19.125 5.52 19.125 5.52 18.955 5.43 18.955 5.43 18.185 2.665 18.185 2.665 17.665 0.085 17.665 0.085 18.955 0 18.955 0 19.125 0.085 19.125 0.085 20.415 ;
      POLYGON 5.43 18.015 5.43 16.405 5.52 16.405 5.52 16.235 5.43 16.235 5.43 14.625 2.835 14.625 2.835 15.145 0.085 15.145 0.085 16.235 0 16.235 0 16.405 0.085 16.405 0.085 17.495 2.835 17.495 2.835 18.015 ;
      RECT 139.38 16.235 139.84 16.405 ;
      POLYGON 2.665 14.975 2.665 14.455 5.43 14.455 5.43 13.685 5.52 13.685 5.52 13.515 3.595 13.515 3.595 12.745 1.735 12.745 1.735 12.225 0.085 12.225 0.085 13.515 0 13.515 0 13.685 0.085 13.685 0.085 14.975 ;
      RECT 139.38 13.515 139.84 13.685 ;
      POLYGON 3.595 12.575 3.595 10.965 3.68 10.965 3.68 10.795 2.675 10.795 2.675 9.185 1.465 9.185 1.465 9.705 0.085 9.705 0.085 10.795 0 10.795 0 10.965 0.085 10.965 0.085 12.055 1.905 12.055 1.905 12.575 ;
      RECT 139.38 10.795 139.84 10.965 ;
      POLYGON 1.295 9.535 1.295 9.015 2.675 9.015 2.675 8.245 2.76 8.245 2.76 8.075 2.675 8.075 2.675 7.305 1.295 7.305 1.295 6.785 0.085 6.785 0.085 8.075 0 8.075 0 8.245 0.085 8.245 0.085 9.535 ;
      RECT 139.38 8.075 139.84 8.245 ;
      POLYGON 2.675 7.135 2.675 5.525 5.52 5.525 5.52 5.355 5.43 5.355 5.43 3.745 2.835 3.745 2.835 4.265 0.085 4.265 0.085 5.355 0 5.355 0 5.525 0.085 5.525 0.085 6.615 1.465 6.615 1.465 7.135 ;
      RECT 139.38 5.355 139.84 5.525 ;
      POLYGON 2.665 4.095 2.665 3.575 5.43 3.575 5.43 2.805 5.52 2.805 5.52 2.635 5.43 2.635 5.43 1.865 2.665 1.865 2.665 1.345 0.085 1.345 0.085 2.635 0 2.635 0 2.805 0.085 2.805 0.085 4.095 ;
      RECT 139.38 2.635 139.84 2.805 ;
      POLYGON 135.155 1.715 135.155 0.085 135.325 0.085 135.325 1.25 135.615 1.25 135.615 0.085 135.785 0.085 135.785 1.175 137.605 1.175 137.605 1.695 139.295 1.695 139.295 0.085 139.84 0.085 139.84 -0.085 0 -0.085 0 0.085 0.085 0.085 0.085 1.175 2.835 1.175 2.835 1.695 5.43 1.695 5.43 0.085 5.605 0.085 5.605 1.175 7.425 1.175 7.425 1.695 9.115 1.695 9.115 0.085 10.205 0.085 10.205 1.25 10.495 1.25 10.495 0.085 10.665 0.085 10.665 1.175 13.415 1.175 13.415 1.695 16.01 1.695 16.01 0.085 16.185 0.085 16.185 1.175 18.935 1.175 18.935 1.695 21.53 1.695 21.53 0.085 21.705 0.085 21.705 1.175 23.085 1.175 23.085 1.695 24.295 1.695 24.295 0.085 24.925 0.085 24.925 1.25 25.215 1.25 25.215 0.085 25.385 0.085 25.385 1.175 28.135 1.175 28.135 1.695 30.73 1.695 30.73 0.085 30.905 0.085 30.905 1.175 33.655 1.175 33.655 1.695 36.25 1.695 36.25 0.085 36.425 0.085 36.425 1.175 37.805 1.175 37.805 1.695 39.015 1.695 39.015 0.085 39.645 0.085 39.645 1.25 39.935 1.25 39.935 0.085 40.105 0.085 40.105 1.175 42.855 1.175 42.855 1.695 45.45 1.695 45.45 0.085 45.625 0.085 45.625 1.175 48.375 1.175 48.375 1.695 50.97 1.695 50.97 0.085 51.145 0.085 51.145 1.175 52.525 1.175 52.525 1.695 53.735 1.695 53.735 0.085 54.365 0.085 54.365 1.25 54.655 1.25 54.655 0.085 54.825 0.085 54.825 1.175 57.575 1.175 57.575 1.695 60.17 1.695 60.17 0.085 60.345 0.085 60.345 1.175 63.095 1.175 63.095 1.695 65.69 1.695 65.69 0.085 65.865 0.085 65.865 1.175 67.245 1.175 67.245 1.695 68.455 1.695 68.455 0.085 69.085 0.085 69.085 1.25 69.375 1.25 69.375 0.085 69.545 0.085 69.545 1.175 72.295 1.175 72.295 1.695 74.89 1.695 74.89 0.085 75.065 0.085 75.065 1.175 77.815 1.175 77.815 1.695 80.41 1.695 80.41 0.085 80.585 0.085 80.585 1.175 81.965 1.175 81.965 1.695 83.175 1.695 83.175 0.085 83.805 0.085 83.805 1.25 84.095 1.25 84.095 0.085 85.155 0.085 85.155 0.585 85.485 0.585 85.485 0.085 86.49 0.085 86.49 0.545 86.74 0.545 86.74 0.085 88.63 0.085 88.63 0.515 88.96 0.515 88.96 0.085 89.595 0.085 89.595 0.545 89.965 0.545 89.965 0.085 91.58 0.085 91.58 0.545 91.83 0.545 91.83 0.085 92.35 0.085 92.35 0.465 92.68 0.465 92.68 0.085 93.02 0.085 93.02 1.225 93.325 1.225 93.325 0.085 93.925 0.085 93.925 1.175 95.745 1.175 95.745 1.695 97.435 1.695 97.435 0.085 98.525 0.085 98.525 1.25 98.815 1.25 98.815 0.085 98.985 0.085 98.985 1.175 101.735 1.175 101.735 1.695 104.33 1.695 104.33 0.085 104.505 0.085 104.505 1.175 107.255 1.175 107.255 1.695 109.85 1.695 109.85 0.085 110.025 0.085 110.025 1.175 111.405 1.175 111.405 1.695 112.615 1.695 112.615 0.085 113.245 0.085 113.245 1.25 113.535 1.25 113.535 0.085 113.705 0.085 113.705 1.175 116.455 1.175 116.455 1.695 119.05 1.695 119.05 0.085 119.225 0.085 119.225 1.175 121.975 1.175 121.975 1.695 124.57 1.695 124.57 0.085 124.745 0.085 124.745 1.175 126.125 1.175 126.125 1.695 127.335 1.695 127.335 0.085 127.965 0.085 127.965 1.25 128.255 1.25 128.255 0.085 128.425 0.085 128.425 1.175 131.175 1.175 131.175 1.695 133.77 1.695 133.77 0.085 133.945 0.085 133.945 1.175 134.635 1.175 134.635 1.715 ;
      POLYGON 108.39 103.19 108.39 86.87 139.67 86.87 139.67 0.17 0.17 0.17 0.17 86.87 31.45 86.87 31.45 103.19 ;
    LAYER via ;
      RECT 103.365 103.165 103.515 103.315 ;
      RECT 103.045 103.165 103.195 103.315 ;
      RECT 102.725 103.165 102.875 103.315 ;
      RECT 102.405 103.165 102.555 103.315 ;
      RECT 72.125 103.165 72.275 103.315 ;
      RECT 71.805 103.165 71.955 103.315 ;
      RECT 71.485 103.165 71.635 103.315 ;
      RECT 71.165 103.165 71.315 103.315 ;
      RECT 40.885 103.165 41.035 103.315 ;
      RECT 40.565 103.165 40.715 103.315 ;
      RECT 40.245 103.165 40.395 103.315 ;
      RECT 39.925 103.165 40.075 103.315 ;
      RECT 75.295 102.535 75.445 102.685 ;
      RECT 73.295 102.535 73.445 102.685 ;
      RECT 68.695 102.195 68.845 102.345 ;
      RECT 127.365 86.845 127.515 86.995 ;
      RECT 127.045 86.845 127.195 86.995 ;
      RECT 126.725 86.845 126.875 86.995 ;
      RECT 126.405 86.845 126.555 86.995 ;
      RECT 20.485 86.845 20.635 86.995 ;
      RECT 20.165 86.845 20.315 86.995 ;
      RECT 19.845 86.845 19.995 86.995 ;
      RECT 19.525 86.845 19.675 86.995 ;
      RECT 139.525 78.805 139.675 78.955 ;
      RECT 0.165 78.805 0.315 78.955 ;
      RECT 139.525 54.505 139.675 54.655 ;
      RECT 0.165 54.505 0.315 54.655 ;
      RECT 139.525 35.285 139.675 35.435 ;
      RECT 0.165 35.285 0.315 35.435 ;
      RECT 139.525 10.805 139.675 10.955 ;
      RECT 0.165 10.805 0.315 10.955 ;
      RECT 66.395 1.555 66.545 1.705 ;
      RECT 127.365 0.045 127.515 0.195 ;
      RECT 127.045 0.045 127.195 0.195 ;
      RECT 126.725 0.045 126.875 0.195 ;
      RECT 126.405 0.045 126.555 0.195 ;
      RECT 103.365 0.045 103.515 0.195 ;
      RECT 103.045 0.045 103.195 0.195 ;
      RECT 102.725 0.045 102.875 0.195 ;
      RECT 102.405 0.045 102.555 0.195 ;
      RECT 72.125 0.045 72.275 0.195 ;
      RECT 71.805 0.045 71.955 0.195 ;
      RECT 71.485 0.045 71.635 0.195 ;
      RECT 71.165 0.045 71.315 0.195 ;
      RECT 40.885 0.045 41.035 0.195 ;
      RECT 40.565 0.045 40.715 0.195 ;
      RECT 40.245 0.045 40.395 0.195 ;
      RECT 39.925 0.045 40.075 0.195 ;
      RECT 20.485 0.045 20.635 0.195 ;
      RECT 20.165 0.045 20.315 0.195 ;
      RECT 19.845 0.045 19.995 0.195 ;
      RECT 19.525 0.045 19.675 0.195 ;
    LAYER via2 ;
      RECT 103.26 103.14 103.46 103.34 ;
      RECT 102.86 103.14 103.06 103.34 ;
      RECT 102.46 103.14 102.66 103.34 ;
      RECT 72.02 103.14 72.22 103.34 ;
      RECT 71.62 103.14 71.82 103.34 ;
      RECT 71.22 103.14 71.42 103.34 ;
      RECT 40.78 103.14 40.98 103.34 ;
      RECT 40.38 103.14 40.58 103.34 ;
      RECT 39.98 103.14 40.18 103.34 ;
      RECT 101.33 102.43 101.53 102.63 ;
      RECT 69.59 102.43 69.79 102.63 ;
      RECT 34.63 101.9 34.83 102.1 ;
      RECT 92.29 101.75 92.49 101.95 ;
      RECT 63.77 101.75 63.97 101.95 ;
      RECT 43.07 101.75 43.27 101.95 ;
      RECT 127.26 86.82 127.46 87.02 ;
      RECT 126.86 86.82 127.06 87.02 ;
      RECT 126.46 86.82 126.66 87.02 ;
      RECT 20.38 86.82 20.58 87.02 ;
      RECT 19.98 86.82 20.18 87.02 ;
      RECT 19.58 86.82 19.78 87.02 ;
      RECT 21.29 86.11 21.49 86.31 ;
      RECT 1.28 82.45 1.48 82.65 ;
      RECT 139.5 78.78 139.7 78.98 ;
      RECT 0.14 78.78 0.34 78.98 ;
      RECT 1.28 71.57 1.48 71.77 ;
      RECT 139.5 54.48 139.7 54.68 ;
      RECT 0.14 54.48 0.34 54.68 ;
      RECT 1.28 52.53 1.48 52.73 ;
      RECT 1.28 42.33 1.48 42.53 ;
      RECT 139.5 35.26 139.7 35.46 ;
      RECT 0.14 35.26 0.34 35.46 ;
      RECT 1.28 33.49 1.48 33.69 ;
      RECT 1.67 29.67 1.87 29.87 ;
      RECT 1.28 25.33 1.48 25.53 ;
      RECT 1.28 15.13 1.48 15.33 ;
      RECT 139.5 10.78 139.7 10.98 ;
      RECT 0.14 10.78 0.34 10.98 ;
      RECT 1.28 6.97 1.48 7.17 ;
      RECT 127.26 0.02 127.46 0.22 ;
      RECT 126.86 0.02 127.06 0.22 ;
      RECT 126.46 0.02 126.66 0.22 ;
      RECT 103.26 0.02 103.46 0.22 ;
      RECT 102.86 0.02 103.06 0.22 ;
      RECT 102.46 0.02 102.66 0.22 ;
      RECT 72.02 0.02 72.22 0.22 ;
      RECT 71.62 0.02 71.82 0.22 ;
      RECT 71.22 0.02 71.42 0.22 ;
      RECT 40.78 0.02 40.98 0.22 ;
      RECT 40.38 0.02 40.58 0.22 ;
      RECT 39.98 0.02 40.18 0.22 ;
      RECT 20.38 0.02 20.58 0.22 ;
      RECT 19.98 0.02 20.18 0.22 ;
      RECT 19.58 0.02 19.78 0.22 ;
    LAYER via3 ;
      RECT 103.26 103.14 103.46 103.34 ;
      RECT 102.86 103.14 103.06 103.34 ;
      RECT 102.46 103.14 102.66 103.34 ;
      RECT 72.02 103.14 72.22 103.34 ;
      RECT 71.62 103.14 71.82 103.34 ;
      RECT 71.22 103.14 71.42 103.34 ;
      RECT 40.78 103.14 40.98 103.34 ;
      RECT 40.38 103.14 40.58 103.34 ;
      RECT 39.98 103.14 40.18 103.34 ;
      RECT 93.59 101.75 93.79 101.95 ;
      RECT 51.88 101.75 52.08 101.95 ;
      RECT 127.26 86.82 127.46 87.02 ;
      RECT 126.86 86.82 127.06 87.02 ;
      RECT 126.46 86.82 126.66 87.02 ;
      RECT 20.38 86.82 20.58 87.02 ;
      RECT 19.98 86.82 20.18 87.02 ;
      RECT 19.58 86.82 19.78 87.02 ;
      RECT 139.5 78.78 139.7 78.98 ;
      RECT 0.14 78.78 0.34 78.98 ;
      RECT 139.5 54.48 139.7 54.68 ;
      RECT 0.14 54.48 0.34 54.68 ;
      RECT 139.5 35.26 139.7 35.46 ;
      RECT 0.14 35.26 0.34 35.46 ;
      RECT 1.59 21.51 1.79 21.71 ;
      RECT 139.5 10.78 139.7 10.98 ;
      RECT 0.14 10.78 0.34 10.98 ;
      RECT 127.26 0.02 127.46 0.22 ;
      RECT 126.86 0.02 127.06 0.22 ;
      RECT 126.46 0.02 126.66 0.22 ;
      RECT 103.26 0.02 103.46 0.22 ;
      RECT 102.86 0.02 103.06 0.22 ;
      RECT 102.46 0.02 102.66 0.22 ;
      RECT 72.02 0.02 72.22 0.22 ;
      RECT 71.62 0.02 71.82 0.22 ;
      RECT 71.22 0.02 71.42 0.22 ;
      RECT 40.78 0.02 40.98 0.22 ;
      RECT 40.38 0.02 40.58 0.22 ;
      RECT 39.98 0.02 40.18 0.22 ;
      RECT 20.38 0.02 20.58 0.22 ;
      RECT 19.98 0.02 20.18 0.22 ;
      RECT 19.58 0.02 19.78 0.22 ;
    LAYER via4 ;
      RECT 4.06 80.12 4.86 80.92 ;
      RECT 4.06 78.52 4.86 79.32 ;
      RECT 139.2 78.48 140 79.28 ;
      RECT -0.16 78.48 0.64 79.28 ;
      RECT 4.06 76.92 4.86 77.72 ;
      RECT 139.2 54.18 140 54.98 ;
      RECT -0.16 54.18 0.64 54.98 ;
      RECT 4.06 36.12 4.86 36.92 ;
      RECT 139.2 34.96 140 35.76 ;
      RECT -0.16 34.96 0.64 35.76 ;
      RECT 4.06 34.52 4.86 35.32 ;
      RECT 4.06 32.92 4.86 33.72 ;
      RECT 139.2 10.48 140 11.28 ;
      RECT -0.16 10.48 0.64 11.28 ;
    LAYER OVERLAP ;
      POLYGON 0 0 0 87.04 31.28 87.04 31.28 103.36 108.56 103.36 108.56 87.04 139.84 87.04 139.84 0 ;
  END
END sb_1__0_

END LIBRARY
